`ifndef MACROS_SVH_
`define MACROS_SVH_

`define ADD 5'b0
`define SUB 5'b1
`define XOR 5'b10
`define OR 5'b11
`define AND 5'b100
`define SLL 5'b101
`define SRL 5'b110
`define SRA 5'b111
`define SLT 5'b1000
`define SLTU 5'b1001
// 
`define ADDI 5'b1010
`define XORI 5'b1011
`define ORI 5'b1100
`define ANDI 5'b1101
`define SLLI 5'b1110
`define SRLI 5'b1111
`define SRAI 5'b10000
`define SLTI 5'b10001
`define SLTIU 5'b10010
//
`define UNUSED_FIELD 5'b11110
`define INVALID_INSTRUCTION 5'b11111

`endif

